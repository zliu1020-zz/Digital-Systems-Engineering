----------------------------------------------------------------------
-- begin uw-generated entity for gate shim 
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use ieee.std_logic_1164.all;
entity myflipflop is
  port (
      i_clock  : in STD_LOGIC
    ; i_d  : in STD_LOGIC
    ; i_ce  : in STD_LOGIC
    ; i_reset  : in STD_LOGIC
    ; i_sel  : in STD_LOGIC
    ; i_d2  : in STD_LOGIC
    ; o_q  : out STD_LOGIC
    ; o_q_a  : out STD_LOGIC
    ; o_q_b  : out STD_LOGIC
    ; o_q_c  : out STD_LOGIC
    ; o_q_d  : out STD_LOGIC
  );
end entity;

----------------------------------------------------------------------
-- begin uw-generated architecture for gate shim
----------------------------------------------------------------------

architecture gate_shim of myflipflop is
  signal VDD, VSS : std_logic; 
begin
  gate : entity work.myflipflop_gate
    port map (
        i_clock => i_clock
      , i_d => i_d
      , i_ce => i_ce
      , i_reset => i_reset
      , i_sel => i_sel
      , i_d2 => i_d2
      , o_q => o_q
      , o_q_a => o_q_a
      , o_q_b => o_q_b
      , o_q_c => o_q_c
      , o_q_d => o_q_d
    );
end architecture;

----------------------------------------------------------------------
-- begin uw-generated entity for gate shim 
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use ieee.std_logic_1164.all;
entity myflipflop is
  port (
      i_clock  : in STD_LOGIC
    ; i_d  : in STD_LOGIC
    ; i_ce  : in STD_LOGIC
    ; i_reset  : in STD_LOGIC
    ; i_sel  : in STD_LOGIC
    ; i_d2  : in STD_LOGIC
    ; o_q  : out STD_LOGIC
    ; o_q_a  : out STD_LOGIC
    ; o_q_b  : out STD_LOGIC
    ; o_q_c  : out STD_LOGIC
    ; o_q_d  : out STD_LOGIC
  );
end entity;

----------------------------------------------------------------------
-- begin uw-generated architecture for gate shim
----------------------------------------------------------------------

architecture gate_shim of myflipflop is
  signal VDD, VSS : std_logic; 
begin
  gate : entity work.myflipflop_gate
    port map (
        i_clock => i_clock
      , i_d => i_d
      , i_ce => i_ce
      , i_reset => i_reset
      , i_sel => i_sel
      , i_d2 => i_d2
      , o_q => o_q
      , o_q_a => o_q_a
      , o_q_b => o_q_b
      , o_q_c => o_q_c
      , o_q_d => o_q_d
    );
end architecture;

----------------------------------------------------------------------
-- begin uw-generated entity for gate shim 
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use ieee.std_logic_1164.all;
entity myflipflop is
  port (
      i_clock  : in STD_LOGIC
    ; i_d  : in STD_LOGIC
    ; i_ce  : in STD_LOGIC
    ; i_reset  : in STD_LOGIC
    ; i_sel  : in STD_LOGIC
    ; i_d2  : in STD_LOGIC
    ; o_q  : out STD_LOGIC
    ; o_q_a  : out STD_LOGIC
    ; o_q_b  : out STD_LOGIC
    ; o_q_c  : out STD_LOGIC
    ; o_q_d  : out STD_LOGIC
  );
end entity;

----------------------------------------------------------------------
-- begin uw-generated architecture for gate shim
----------------------------------------------------------------------

architecture gate_shim of myflipflop is
  signal VDD, VSS : std_logic; 
begin
  gate : entity work.myflipflop_gate
    port map (
        i_clock => i_clock
      , i_d => i_d
      , i_ce => i_ce
      , i_reset => i_reset
      , i_sel => i_sel
      , i_d2 => i_d2
      , o_q => o_q
      , o_q_a => o_q_a
      , o_q_b => o_q_b
      , o_q_c => o_q_c
      , o_q_d => o_q_d
    );
end architecture;

----------------------------------------------------------------------
-- begin uw-generated entity for gate shim 
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use ieee.std_logic_1164.all;
entity myflipflop is
  port (
      i_clock  : in STD_LOGIC
    ; i_d  : in STD_LOGIC
    ; i_ce  : in STD_LOGIC
    ; i_reset  : in STD_LOGIC
    ; i_sel  : in STD_LOGIC
    ; i_d2  : in STD_LOGIC
    ; o_q  : out STD_LOGIC
    ; o_q_a  : out STD_LOGIC
    ; o_q_b  : out STD_LOGIC
    ; o_q_c  : out STD_LOGIC
    ; o_q_d  : out STD_LOGIC
  );
end entity;

----------------------------------------------------------------------
-- begin uw-generated architecture for gate shim
----------------------------------------------------------------------

architecture gate_shim of myflipflop is
  signal VDD, VSS : std_logic; 
begin
  gate : entity work.myflipflop_gate
    port map (
        i_clock => i_clock
      , i_d => i_d
      , i_ce => i_ce
      , i_reset => i_reset
      , i_sel => i_sel
      , i_d2 => i_d2
      , o_q => o_q
      , o_q_a => o_q_a
      , o_q_b => o_q_b
      , o_q_c => o_q_c
      , o_q_d => o_q_d
    );
end architecture;

